----------------------------------------------------------------------------------
-- Company: KUL - Group T - RDMA Team
-- Engineer: Tolga Kuntman <kuntmantolga@gmail.com>
-- 
-- Create Date: 22/11/2025 12:09:11 PM
-- Design Name: 
-- Module Name: data_mover_controller_axis_master
-- Project Name: RDMA
-- Target Devices: Kria KR260
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
`timescale 1 ns / 1 ps

	module data_mover_controller_master_stream_v1_0_M00_AXIS #
	(
		// Users to add parameters here

		// User parameters ends
		// Do not modify the parameters beyond this line

		// Width of S_AXIS address bus. The slave accepts the read and write addresses of width C_M_AXIS_TDATA_WIDTH.
		parameter integer C_M_AXIS_TDATA_WIDTH	= 32,
		// Start count is the number of clock cycles the master will wait before initiating/issuing any transaction.
		parameter integer C_M_START_COUNT	= 32
	)
	(
		// Users to add ports here
		input wire start,
		input wire [C_M_AXIS_TDATA_WIDTH-1:0] input_data_0,
		input wire [C_M_AXIS_TDATA_WIDTH-1:0] input_data_1,
		input wire [C_M_AXIS_TDATA_WIDTH-1:0] input_data_2,
		input wire [C_M_AXIS_TDATA_WIDTH-1:0] input_data_3,
		input wire [C_M_AXIS_TDATA_WIDTH-1:0] input_data_4,
		input wire [C_M_AXIS_TDATA_WIDTH-1:0] input_data_5,
		input wire [C_M_AXIS_TDATA_WIDTH-1:0] input_data_6,
		input wire [C_M_AXIS_TDATA_WIDTH-1:0] input_data_7,
		output wire busy,
		// User ports ends
		// Do not modify the ports beyond this line

		// Global ports
		input wire  M_AXIS_ACLK,
		// 
		input wire  M_AXIS_ARESETN,
		// Master Stream Ports. TVALID indicates that the master is driving a valid transfer, A transfer takes place when both TVALID and TREADY are asserted. 
		output wire  M_AXIS_TVALID,
		// TDATA is the primary payload that is used to provide the data that is passing across the interface from the master.
		output wire [C_M_AXIS_TDATA_WIDTH-1 : 0] M_AXIS_TDATA,
		// TSTRB is the byte qualifier that indicates whether the content of the associated byte of TDATA is processed as a data byte or a position byte.
		output wire [(C_M_AXIS_TDATA_WIDTH/8)-1 : 0] M_AXIS_TSTRB,
		// TLAST indicates the boundary of a packet.
		output wire  M_AXIS_TLAST,
		// TREADY indicates that the slave can accept a transfer in the current cycle.
		input wire  M_AXIS_TREADY
	);
	// Total number of output data                                                 
	localparam NUMBER_OF_OUTPUT_WORDS = 8;                                               
	                                                                                     
	// function called clogb2 that returns an integer which has the                      
	// value of the ceiling of the log base 2.                                           
	function integer clogb2 (input integer bit_depth);                                   
	  begin                                                                              
	    for(clogb2=0; bit_depth>0; clogb2=clogb2+1)                                      
	      bit_depth = bit_depth >> 1;                                                    
	  end                                                                                
	endfunction                                                                          
	                                                                                     
	// WAIT_COUNT_BITS is the width of the wait counter.                                 
	localparam integer WAIT_COUNT_BITS = clogb2(C_M_START_COUNT-1);                      
	                                                                                     
	// bit_num gives the minimum number of bits needed to address 'depth' size of FIFO.  
	localparam bit_num  = clogb2(NUMBER_OF_OUTPUT_WORDS);                                
	                                                                                     
	// Define the states of state machine                                                
	// The control state machine oversees the writing of input streaming data to the FIFO,
	// and outputs the streaming data from the FIFO                                      
	parameter [1:0] IDLE = 2'b00,        // This is the initial/idle state, waits for start
	                SEND_STREAM   = 2'b01; // In this state the stream data is output through M_AXIS_TDATA
	                                                                                     
	// State variable                                                                    
	reg [1:0] mst_exec_state;                                                            
	// Example design FIFO read pointer                                                  
	reg [bit_num-1:0] read_pointer;                                                      

	// AXI Stream internal signals
	//wait counter. The master waits for the user defined number of clock cycles before initiating a transfer.
	reg [WAIT_COUNT_BITS-1 : 0] 	count;
	//streaming data valid
	wire  	axis_tvalid;
	//streaming data valid delayed by one clock cycle
	reg  	axis_tvalid_delay;
	//Last of the streaming data 
	wire  	axis_tlast;
	//Last of the streaming data delayed by one clock cycle
	reg  	axis_tlast_delay;
	//FIFO implementation signals
	reg [C_M_AXIS_TDATA_WIDTH-1 : 0] 	stream_data_out;
	wire  	tx_en;
	//The master has issued all the streaming data stored in FIFO
	reg  	tx_done;


	// I/O Connections assignments

	assign M_AXIS_TVALID	= axis_tvalid_delay;
	assign M_AXIS_TDATA	= stream_data_out;
	assign M_AXIS_TLAST	= axis_tlast_delay;
	assign M_AXIS_TSTRB	= {(C_M_AXIS_TDATA_WIDTH/8){1'b1}};


	// Control state machine implementation                             
	always @(posedge M_AXIS_ACLK)                                             
	begin                                                                     
	  if (!M_AXIS_ARESETN)                                                    
	  // Synchronous reset (active low)                                       
	    begin                                                                 
	      mst_exec_state <= IDLE;                                             
	    end                                                                   
	  else                                                                    
	    case (mst_exec_state)                                                 
	      IDLE:                                                               
	        // Wait for start signal to begin transmission
	        if (start)                                                        
	          begin                                                           
	            mst_exec_state <= SEND_STREAM;                                
	          end                                                             
	                                                                          
	      SEND_STREAM:                                                        
	        // Send data until all words transmitted
	        if (tx_done)                                                      
	          begin                                                           
	            mst_exec_state <= IDLE;                                       
	          end                                                             
	    endcase                                                               
	end                                                                       

	// Busy signal indicates transmission in progress
	assign busy = (mst_exec_state == SEND_STREAM);                                                                       


	//tvalid generation
	//axis_tvalid is asserted when the control state machine's state is SEND_STREAM and
	//number of output streaming data is less than the NUMBER_OF_OUTPUT_WORDS.
	assign axis_tvalid = ((mst_exec_state == SEND_STREAM) && (read_pointer < NUMBER_OF_OUTPUT_WORDS));
	                                                                                               
	// AXI tlast generation                                                                        
	// axis_tlast is asserted number of output streaming data is NUMBER_OF_OUTPUT_WORDS-1          
	// (0 to NUMBER_OF_OUTPUT_WORDS-1)                                                             
	assign axis_tlast = (read_pointer == NUMBER_OF_OUTPUT_WORDS-1);                                
	                                                                                               
	                                                                                               
	// Delay the axis_tvalid and axis_tlast signal by one clock cycle                              
	// to match the latency of M_AXIS_TDATA                                                        
	always @(posedge M_AXIS_ACLK)                                                                  
	begin                                                                                          
	  if (!M_AXIS_ARESETN)                                                                         
	    begin                                                                                      
	      axis_tvalid_delay <= 1'b0;                                                               
	      axis_tlast_delay <= 1'b0;                                                                
	    end                                                                                        
	  else                                                                                         
	    begin                                                                                      
	      axis_tvalid_delay <= axis_tvalid;                                                        
	      axis_tlast_delay <= axis_tlast;                                                          
	    end                                                                                        
	end                                                                                            


	//read_pointer pointer

	always@(posedge M_AXIS_ACLK)                                               
	begin                                                                            
	  if(!M_AXIS_ARESETN)                                                            
	    begin                                                                        
	      read_pointer <= 0;                                                         
	      tx_done <= 1'b0;                                                           
	    end
	  else if (start && mst_exec_state == IDLE)
	    begin
	      // Reset for new transfer
	      read_pointer <= 0;
	      tx_done <= 1'b0;
	    end
	  else                                                                           
	    if (read_pointer <= NUMBER_OF_OUTPUT_WORDS-1)                                
	      begin                                                                      
	        if (tx_en)                                                               
	          // read pointer is incremented after every read from the FIFO          
	          // when FIFO read signal is enabled.                                   
	          begin                                                                  
	            read_pointer <= read_pointer + 1;                                    
	            tx_done <= 1'b0;                                                     
	          end       
			  else																	
	        begin                                                                    
	          read_pointer <= read_pointer;                                          
	          tx_done <= 1'b0;                                                     
	        end                                                             
	      end                                                                        
	    else if (read_pointer == NUMBER_OF_OUTPUT_WORDS)                             
	      begin                                                                      
	        // tx_done is asserted when NUMBER_OF_OUTPUT_WORDS numbers of streaming data
	        // has been out.                                                         
	        tx_done <= 1'b1;                                                         
	      end                                                                        
	end                                                                              


	// Internal data buffer to hold input data
	reg [C_M_AXIS_TDATA_WIDTH-1:0] data_buffer [0:NUMBER_OF_OUTPUT_WORDS-1];

	// Capture input data when start is asserted
	always @(posedge M_AXIS_ACLK)
	begin
	  if (!M_AXIS_ARESETN)
	    begin
	      data_buffer[0] <= 0;
	      data_buffer[1] <= 0;
	      data_buffer[2] <= 0;
	      data_buffer[3] <= 0;
	      data_buffer[4] <= 0;
	      data_buffer[5] <= 0;
	      data_buffer[6] <= 0;
	      data_buffer[7] <= 0;
	    end
	  else if (start && mst_exec_state == IDLE)
	    begin
	      data_buffer[0] <= input_data_0;
	      data_buffer[1] <= input_data_1;
	      data_buffer[2] <= input_data_2;
	      data_buffer[3] <= input_data_3;
	      data_buffer[4] <= input_data_4;
	      data_buffer[5] <= input_data_5;
	      data_buffer[6] <= input_data_6;
	      data_buffer[7] <= input_data_7;
	    end
	end

	//FIFO read enable generation 
	assign tx_en = M_AXIS_TREADY && axis_tvalid;   
	                                                     
	// Streaming output data from buffer
	always @(posedge M_AXIS_ACLK)                  
	begin                                            
	  if(!M_AXIS_ARESETN)                            
	    begin                                        
	      stream_data_out <= 0;                      
	    end                                          
	  else if (tx_en)  
	    begin                                        
	      stream_data_out <= data_buffer[read_pointer];   
	    end                                          
	end                                              

	// Add user logic here

	// User logic ends

	endmodule